module Testbench(

);

endmodule
