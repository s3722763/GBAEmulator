module Ander (
    input A,
    input B,
    output var C
);
    assign C = A & B;
endmodule